VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_customcell
  CLASS CORE ;
  FOREIGN sky130_customcell ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SITE unithd ;
  PIN in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 2.265 1.580 2.435 ;
        RECT 0.125 0.990 0.895 1.320 ;
        RECT 0.720 0.515 0.895 0.990 ;
        RECT 1.065 0.515 1.235 2.265 ;
        RECT 0.720 0.345 1.235 0.515 ;
        RECT 1.410 0.515 1.580 2.265 ;
        RECT 1.750 2.265 2.265 2.435 ;
        RECT 1.750 0.515 1.920 2.265 ;
        RECT 1.410 0.345 1.920 0.515 ;
        RECT 2.095 0.515 2.265 2.265 ;
        RECT 2.435 2.265 2.950 2.435 ;
        RECT 2.435 0.515 2.605 2.265 ;
        RECT 2.095 0.345 2.605 0.515 ;
        RECT 2.780 0.515 2.950 2.265 ;
        RECT 3.120 2.265 3.635 2.435 ;
        RECT 3.120 0.515 3.290 2.265 ;
        RECT 2.780 0.345 3.290 0.515 ;
        RECT 3.465 0.515 3.635 2.265 ;
        RECT 4.365 1.250 4.700 1.305 ;
        RECT 3.805 1.080 4.700 1.250 ;
        RECT 3.805 0.515 3.975 1.080 ;
        RECT 3.465 0.345 3.975 0.515 ;
    END
  END in
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.243600 ;
    PORT
      LAYER li1 ;
        RECT 5.860 2.265 6.375 2.435 ;
        RECT 4.870 1.345 5.040 2.140 ;
        RECT 4.870 1.085 5.690 1.345 ;
        RECT 4.870 0.445 5.040 1.085 ;
        RECT 5.520 0.515 5.690 1.085 ;
        RECT 5.860 0.515 6.030 2.265 ;
        RECT 5.520 0.345 6.030 0.515 ;
        RECT 6.205 0.515 6.375 2.265 ;
        RECT 6.545 2.265 7.060 2.435 ;
        RECT 6.545 0.515 6.715 2.265 ;
        RECT 6.205 0.345 6.715 0.515 ;
        RECT 6.890 0.515 7.060 2.265 ;
        RECT 7.230 2.265 7.745 2.435 ;
        RECT 7.230 0.515 7.400 2.265 ;
        RECT 6.890 0.345 7.400 0.515 ;
        RECT 7.575 0.515 7.745 2.265 ;
        RECT 7.915 2.265 8.430 2.435 ;
        RECT 7.915 0.515 8.085 2.265 ;
        RECT 7.575 0.345 8.085 0.515 ;
        RECT 8.260 0.555 8.430 2.265 ;
        RECT 8.660 0.555 8.890 1.290 ;
        RECT 8.260 0.345 8.890 0.555 ;
      LAYER mcon ;
        RECT 4.870 1.760 5.040 2.060 ;
        RECT 4.870 0.525 5.040 0.825 ;
        RECT 8.690 1.100 8.860 1.270 ;
      LAYER met1 ;
        RECT 4.840 1.700 5.070 2.120 ;
        RECT 8.625 0.965 8.920 1.300 ;
        RECT 4.840 0.465 5.070 0.885 ;
    END
  END out
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 4.430 1.680 4.600 2.140 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 4.430 1.760 4.600 2.060 ;
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
        RECT 4.400 1.700 4.630 2.480 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 4.430 0.445 4.600 0.905 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 4.430 0.525 4.600 0.825 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
      LAYER met1 ;
        RECT 4.400 0.240 4.630 0.885 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.235 9.390 2.910 ;
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 -0.085 9.195 1.070 ;
    END
  END VNB
END sky130_customcell
END LIBRARY

