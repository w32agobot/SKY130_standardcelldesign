magic
tech sky130A
magscale 1 2
timestamp 1663107964
<< nwell >>
rect -38 247 1878 582
<< pwell >>
rect 1 -17 1839 214
<< nmos >>
rect 932 93 962 177
<< pmos >>
rect 932 340 962 424
<< ndiff >>
rect 874 165 932 177
rect 874 105 886 165
rect 920 105 932 165
rect 874 93 932 105
rect 962 165 1020 177
rect 962 105 974 165
rect 1008 105 1020 165
rect 962 93 1020 105
<< pdiff >>
rect 874 412 932 424
rect 874 352 886 412
rect 920 352 932 412
rect 874 340 932 352
rect 962 412 1020 424
rect 962 352 974 412
rect 1008 352 1020 412
rect 962 340 1020 352
<< ndiffc >>
rect 886 105 920 165
rect 974 105 1008 165
<< pdiffc >>
rect 886 352 920 412
rect 974 352 1008 412
<< poly >>
rect 932 424 962 450
rect 932 271 962 340
rect 931 269 962 271
rect 25 248 147 264
rect 25 214 35 248
rect 70 214 147 248
rect 873 259 962 269
rect 873 225 890 259
rect 924 225 962 259
rect 873 214 962 225
rect 25 198 147 214
rect 932 177 962 214
rect 932 67 962 93
<< polycont >>
rect 35 214 70 248
rect 890 225 924 259
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 213 453 316 487
rect 25 248 179 264
rect 25 214 35 248
rect 70 214 179 248
rect 25 198 179 214
rect 144 103 179 198
rect 213 103 247 453
rect 144 69 247 103
rect 282 103 316 453
rect 350 453 453 487
rect 350 103 384 453
rect 282 69 384 103
rect 419 103 453 453
rect 487 453 590 487
rect 487 103 521 453
rect 419 69 521 103
rect 556 103 590 453
rect 624 453 727 487
rect 624 103 658 453
rect 556 69 658 103
rect 693 103 727 453
rect 1172 453 1275 487
rect 886 412 920 428
rect 886 336 920 352
rect 974 412 1008 428
rect 974 269 1008 352
rect 873 259 940 261
rect 873 250 890 259
rect 761 225 890 250
rect 924 225 940 259
rect 761 216 940 225
rect 974 217 1138 269
rect 761 103 795 216
rect 693 69 795 103
rect 886 165 920 181
rect 886 89 920 105
rect 974 165 1008 217
rect 974 89 1008 105
rect 1104 103 1138 217
rect 1172 103 1206 453
rect 1104 69 1206 103
rect 1241 103 1275 453
rect 1309 453 1412 487
rect 1309 103 1343 453
rect 1241 69 1343 103
rect 1378 103 1412 453
rect 1446 453 1549 487
rect 1446 103 1480 453
rect 1378 69 1480 103
rect 1515 103 1549 453
rect 1583 453 1686 487
rect 1583 103 1617 453
rect 1515 69 1617 103
rect 1652 111 1686 453
rect 1732 254 1778 258
rect 1732 220 1738 254
rect 1772 220 1778 254
rect 1732 111 1778 220
rect 1652 69 1778 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 886 352 920 412
rect 974 352 1008 412
rect 886 105 920 165
rect 974 105 1008 165
rect 1738 220 1772 254
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 880 412 926 496
rect 880 352 886 412
rect 920 352 926 412
rect 880 340 926 352
rect 968 412 1014 424
rect 968 352 974 412
rect 1008 352 1014 412
rect 968 340 1014 352
rect 1725 254 1784 260
rect 1725 220 1738 254
rect 1772 220 1784 254
rect 1725 193 1784 220
rect 880 165 926 177
rect 880 105 886 165
rect 920 105 926 165
rect 880 48 926 105
rect 968 165 1014 177
rect 968 105 974 165
rect 1008 105 1014 165
rect 968 93 1014 105
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel metal1 s 0 496 1840 592 0 FreeSans 160 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 213 527 247 561 0 FreeSans 160 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 213 -17 247 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 0 -48 1840 48 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 213 527 247 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 213 -17 247 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 1738 220 1772 254 0 FreeSans 160 0 0 0 out
port 2 nsew signal output
flabel locali s 38 221 72 255 7 FreeSans 160 0 0 0 in
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1840 544
string LEFclass CORE
string LEForigin 0 0
string LEFsite unithd
string LEFsource USER
<< end >>
